module R4Booth #(
    parameter PARM_MANT = 23 // Width of the mantissa
) (
    input [PARM_MANT : 0] MantA_i, // Input multiplicand (24 bits: hidden bit + mantissa)
    input [PARM_MANT : 0] MantB_i, // Input multiplier (24 bits: hidden bit + mantissa)

    output [2*PARM_MANT + 2 : 0] pp_00_o, // Partial product outputs (49 bits each)
    output [2*PARM_MANT + 2 : 0] pp_01_o,
    output [2*PARM_MANT + 2 : 0] pp_02_o,
    output [2*PARM_MANT + 2 : 0] pp_03_o,
    output [2*PARM_MANT + 2 : 0] pp_04_o,
    output [2*PARM_MANT + 2 : 0] pp_05_o,
    output [2*PARM_MANT + 2 : 0] pp_06_o,
    output [2*PARM_MANT + 2 : 0] pp_07_o,
    output [2*PARM_MANT + 2 : 0] pp_08_o,
    output [2*PARM_MANT + 2 : 0] pp_09_o,
    output [2*PARM_MANT + 2 : 0] pp_10_o,
    output [2*PARM_MANT + 2 : 0] pp_11_o,
    output [2*PARM_MANT + 1 : 0] pp_12_o
);

    // Number of partial products generated by Booth's algorithm
    parameter PARM_PP = ((PARM_MANT + 1) + 1 + 1) / 2;

    // Extend the multiplier with padding for Booth encoding
    wire [PARM_MANT + 3 : 0] mant_B_Padding = {2'd0, MantB_i, 1'd0};

    // Booth encoding signals
    wire [PARM_PP - 1 : 0] mul1x;    // Indicates a 1x multiplicand
    wire [PARM_PP - 1 : 0] mul2x;    // Indicates a 2x multiplicand
    wire [PARM_PP - 1 : 0] mulsign;  // Indicates a negative multiplicand

    // Generate Booth encoding for each partial product
    generate
        genvar j;
        for (j = 0; j < 13; j = j + 1) begin
            assign mul1x[j] = mant_B_Padding[j*2] ^ mant_B_Padding[j*2 + 1]; // XOR for 1x
            assign mul2x[j] = ((~mant_B_Padding[j*2]) & (~mant_B_Padding[j*2 + 1]) & mant_B_Padding[j*2 + 2]) ||
                              (mant_B_Padding[j*2] & mant_B_Padding[j*2 + 1] & ~mant_B_Padding[j*2 + 2]); // Detect 2x
            assign mulsign[j] = mant_B_Padding[j*2 + 2]; // Sign bit
        end
    endgenerate

    // Temporary storage for partial products
    reg [PARM_MANT + 1 : 0] booth_PP_tmp [PARM_PP - 1 : 0];
    wire [PARM_MANT + 1 : 0] booth_PP [PARM_PP - 1 : 0];

    // Generate partial products based on Booth encoding
    integer idx;
    always @(*) begin
        for (idx = 0; idx < PARM_PP; idx = idx + 1) begin
            if (mul1x[idx]) 
                booth_PP_tmp[idx] = MantA_i; // 1x multiplicand
            else if (mul2x[idx]) 
                booth_PP_tmp[idx] = MantA_i << 1; // 2x multiplicand
            else 
                booth_PP_tmp[idx] = 0; // No multiplicand
        end
    end

    // Apply sign correction to partial products (2's complement for negative values)
    generate
        genvar k;
        for (k = 0; k < PARM_PP; k = k + 1) begin
            assign booth_PP[k] = (mulsign[k]) ? ~booth_PP_tmp[k] : booth_PP_tmp[k];
        end
    endgenerate

    // Generate final partial products with proper alignment
    assign pp_00_o = {21'd0, ~mulsign[0], {2{mulsign[0]}}, booth_PP[0]};
    assign pp_01_o = {21'd1, ~mulsign[1], booth_PP[1], 1'b0, mulsign[0]};
    assign pp_02_o = {19'd1, ~mulsign[2], booth_PP[2], 1'b0, mulsign[1], 2'd0};
    assign pp_03_o = {17'd1, ~mulsign[3], booth_PP[3], 1'b0, mulsign[2], 4'd0};
    assign pp_04_o = {15'd1, ~mulsign[4], booth_PP[4], 1'b0, mulsign[3], 6'd0};
    assign pp_05_o = {13'd1, ~mulsign[5], booth_PP[5], 1'b0, mulsign[4], 8'd0};
    assign pp_06_o = {11'd1, ~mulsign[6], booth_PP[6], 1'b0, mulsign[5], 10'd0};
    assign pp_07_o = {9'd1, ~mulsign[7], booth_PP[7], 1'b0, mulsign[6], 12'd0};
    assign pp_08_o = {7'd1, ~mulsign[8], booth_PP[8], 1'b0, mulsign[7], 14'd0};
    assign pp_09_o = {5'd1, ~mulsign[9], booth_PP[9], 1'b0, mulsign[8], 16'd0};
    assign pp_10_o = {3'd1, ~mulsign[10], booth_PP[10], 1'b0, mulsign[9], 18'd0};
    assign pp_11_o = {1'd1, ~mulsign[11], booth_PP[11], 1'b0, mulsign[10], 20'd0};
    assign pp_12_o = {booth_PP[12][PARM_MANT : 0], 1'b0, mulsign[11], 22'd0}; // Save one bit, MSB is always 0

endmodule
