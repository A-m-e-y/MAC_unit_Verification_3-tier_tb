module tb;

initial begin
    // Testbench code goes here
    $display("Testbench started");
    
    // Add your test cases and verification logic here
    
    // End of testbench
    $display("Testbench completed");
    $finish;    
end

endmodule